module complex_multiplier(
	input           clk, // input clk
	input   [15:0]  ar,  // input [15 : 0] ar
	input   [15:0]  ai,  // input [15 : 0] ai
	input   [15:0]  br,  // input [15 : 0] br
	input   [15:0]  bi,  // input [15 : 0] bi
	output  [32:0]  pr,  // output [32 : 0] pr
	output  [32:0]  pi   // output [32 : 0] pi

); 
endmodule
